
module tcm_mem_ram
(
    // Inputs
     input           clk0_i
    ,input           rst0_i
    ,input  [ 13:0]  addr0_i
    ,input  [ 31:0]  data0_i
    ,input  [  3:0]  wr0_i
    ,input           clk1_i
    ,input           rst1_i
    ,input  [ 13:0]  addr1_i
    ,input  [ 31:0]  data1_i
    ,input  [  3:0]  wr1_i

    // Outputs
    ,output [ 31:0]  data0_o
    ,output [ 31:0]  data1_o
);



//-----------------------------------------------------------------
// Dual Port RAM 64KB
// Mode: Read First
//-----------------------------------------------------------------
/* verilator lint_off MULTIDRIVEN */
localparam MEMSIZE = 32;
reg [31:0]   ram [0:MEMSIZE-1] /*verilator public*/;
/* verilator lint_on MULTIDRIVEN */

reg [31:0] ram_read0_q;
reg [31:0] ram_read1_q;

// Synchronous write
always @ (posedge clk0_i)
begin
    if (rst0_i) ;
    else begin

        if (addr0_i < MEMSIZE*4)
        begin
            if (wr0_i[0])
                ram[addr0_i][7:0] <= data0_i[7:0];
            if (wr0_i[1])
                ram[addr0_i][15:8] <= data0_i[15:8];
            if (wr0_i[2])
                ram[addr0_i][23:16] <= data0_i[23:16];
            if (wr0_i[3])
                ram[addr0_i][31:24] <= data0_i[31:24];
            ram_read0_q <= ram[addr0_i];
        end else ram_read0_q <= 32'd0;
        
        if (addr1_i < MEMSIZE*4)
        begin
            if (wr1_i[0])
                ram[addr1_i][7:0] <= data1_i[7:0];
            if (wr1_i[1])
                ram[addr1_i][15:8] <= data1_i[15:8];
            if (wr1_i[2])
                ram[addr1_i][23:16] <= data1_i[23:16];
            if (wr1_i[3])
                ram[addr1_i][31:24] <= data1_i[31:24];
            ram_read1_q <= ram[addr1_i];
        end else ram_read1_q <= 32'd0;
    end
end

assign data0_o = ram_read0_q;
assign data1_o = ram_read1_q;



endmodule
